library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity anode_switcher is
    Port ( clock : in  STD_LOGIC;
           reset : in  STD_LOGIC;
           enable : in  STD_LOGIC;
           anode : out  STD_LOGIC_VECTOR (3 downto 0));
end anode_switcher;

architecture Behavioral of anode_switcher is
begin
		


end Behavioral;

